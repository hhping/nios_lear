// kernel.v

// Generated using ACDS version 14.1 186 at 2018.08.23.22:26:26

`timescale 1 ps / 1 ps
module kernel (
		input  wire        clk_clk,          //        clk.clk
		output wire        epcs_flash_dclk,  // epcs_flash.dclk
		output wire        epcs_flash_sce,   //           .sce
		output wire        epcs_flash_sdo,   //           .sdo
		input  wire        epcs_flash_data0, //           .data0
		input  wire        reset_reset_n,    //      reset.reset_n
		output wire [13:0] sdram_ctrl_addr,  // sdram_ctrl.addr
		output wire [1:0]  sdram_ctrl_ba,    //           .ba
		output wire        sdram_ctrl_cas_n, //           .cas_n
		output wire        sdram_ctrl_cke,   //           .cke
		output wire        sdram_ctrl_cs_n,  //           .cs_n
		inout  wire [15:0] sdram_ctrl_dq,    //           .dq
		output wire [1:0]  sdram_ctrl_dqm,   //           .dqm
		output wire        sdram_ctrl_ras_n, //           .ras_n
		output wire        sdram_ctrl_we_n,  //           .we_n
		input  wire        uart_rxd,         //       uart.rxd
		output wire        uart_txd          //           .txd
	);

	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [27:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                             // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_0_cf_0_ctl_chipselect;                     // mm_interconnect_0:cf_0_ctl_chipselect -> cf_0:av_ctl_chipselect_n
	wire   [3:0] mm_interconnect_0_cf_0_ctl_readdata;                       // cf_0:av_ctl_readdata -> mm_interconnect_0:cf_0_ctl_readdata
	wire   [1:0] mm_interconnect_0_cf_0_ctl_address;                        // mm_interconnect_0:cf_0_ctl_address -> cf_0:av_ctl_address
	wire         mm_interconnect_0_cf_0_ctl_read;                           // mm_interconnect_0:cf_0_ctl_read -> cf_0:av_ctl_read_n
	wire         mm_interconnect_0_cf_0_ctl_write;                          // mm_interconnect_0:cf_0_ctl_write -> cf_0:av_ctl_write_n
	wire   [3:0] mm_interconnect_0_cf_0_ctl_writedata;                      // mm_interconnect_0:cf_0_ctl_writedata -> cf_0:av_ctl_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_epcs_epcs_control_port_chipselect;       // mm_interconnect_0:epcs_epcs_control_port_chipselect -> epcs:chipselect
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_readdata;         // epcs:readdata -> mm_interconnect_0:epcs_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_epcs_control_port_address;          // mm_interconnect_0:epcs_epcs_control_port_address -> epcs:address
	wire         mm_interconnect_0_epcs_epcs_control_port_read;             // mm_interconnect_0:epcs_epcs_control_port_read -> epcs:read_n
	wire         mm_interconnect_0_epcs_epcs_control_port_write;            // mm_interconnect_0:epcs_epcs_control_port_write -> epcs:write_n
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_writedata;        // mm_interconnect_0:epcs_epcs_control_port_writedata -> epcs:writedata
	wire         mm_interconnect_0_cf_0_ide_chipselect;                     // mm_interconnect_0:cf_0_ide_chipselect -> cf_0:av_ide_chipselect_n
	wire  [15:0] mm_interconnect_0_cf_0_ide_readdata;                       // cf_0:av_ide_readdata -> mm_interconnect_0:cf_0_ide_readdata
	wire   [3:0] mm_interconnect_0_cf_0_ide_address;                        // mm_interconnect_0:cf_0_ide_address -> cf_0:av_ide_address
	wire         mm_interconnect_0_cf_0_ide_read;                           // mm_interconnect_0:cf_0_ide_read -> cf_0:av_ide_read_n
	wire         mm_interconnect_0_cf_0_ide_write;                          // mm_interconnect_0:cf_0_ide_write -> cf_0:av_ide_write_n
	wire  [15:0] mm_interconnect_0_cf_0_ide_writedata;                      // mm_interconnect_0:cf_0_ide_writedata -> cf_0:av_ide_writedata
	wire         mm_interconnect_0_uart_s1_chipselect;                      // mm_interconnect_0:uart_s1_chipselect -> uart:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                        // uart:readdata -> mm_interconnect_0:uart_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                         // mm_interconnect_0:uart_s1_address -> uart:address
	wire         mm_interconnect_0_uart_s1_read;                            // mm_interconnect_0:uart_s1_read -> uart:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;                   // mm_interconnect_0:uart_s1_begintransfer -> uart:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                           // mm_interconnect_0:uart_s1_write -> uart:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                       // mm_interconnect_0:uart_s1_writedata -> uart:writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;             // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;               // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory_s1_address;                // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;             // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                  // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;              // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                  // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_sdram_ctrl_s1_chipselect;                // mm_interconnect_0:sdram_ctrl_s1_chipselect -> sdram_ctrl:az_cs
	wire  [15:0] mm_interconnect_0_sdram_ctrl_s1_readdata;                  // sdram_ctrl:za_data -> mm_interconnect_0:sdram_ctrl_s1_readdata
	wire         mm_interconnect_0_sdram_ctrl_s1_waitrequest;               // sdram_ctrl:za_waitrequest -> mm_interconnect_0:sdram_ctrl_s1_waitrequest
	wire  [25:0] mm_interconnect_0_sdram_ctrl_s1_address;                   // mm_interconnect_0:sdram_ctrl_s1_address -> sdram_ctrl:az_addr
	wire         mm_interconnect_0_sdram_ctrl_s1_read;                      // mm_interconnect_0:sdram_ctrl_s1_read -> sdram_ctrl:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_ctrl_s1_byteenable;                // mm_interconnect_0:sdram_ctrl_s1_byteenable -> sdram_ctrl:az_be_n
	wire         mm_interconnect_0_sdram_ctrl_s1_readdatavalid;             // sdram_ctrl:za_valid -> mm_interconnect_0:sdram_ctrl_s1_readdatavalid
	wire         mm_interconnect_0_sdram_ctrl_s1_write;                     // mm_interconnect_0:sdram_ctrl_s1_write -> sdram_ctrl:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_ctrl_s1_writedata;                 // mm_interconnect_0:sdram_ctrl_s1_writedata -> sdram_ctrl:az_data
	wire         irq_mapper_receiver0_irq;                                  // cf_0:av_ctl_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // cf_0:av_ide_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // uart:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                  // epcs:irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [cf_0:av_reset_n, cpu:reset_n, epcs:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_translator:in_reset, sdram_ctrl:reset_n, sysid:reset_n, uart:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu:reset_req, epcs:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                             // cpu:debug_reset_request -> rst_controller:reset_in1

	kernel_cf_0 cf_0 (
		.clk                 (clk_clk),                                //      clk.clk
		.data_cf             (),                                       // external.export
		.we_n                (),                                       //         .export
		.rfu                 (),                                       //         .export
		.reset_n_cf          (),                                       //         .export
		.power               (),                                       //         .export
		.iowr_n              (),                                       //         .export
		.iord_n              (),                                       //         .export
		.cs_n                (),                                       //         .export
		.addr                (),                                       //         .export
		.iordy               (),                                       //         .export
		.intrq               (),                                       //         .export
		.detect_n            (),                                       //         .export
		.atasel_n            (),                                       //         .export
		.av_reset_n          (~rst_controller_reset_out_reset),        //    reset.reset_n
		.av_ide_chipselect_n (~mm_interconnect_0_cf_0_ide_chipselect), //      ide.chipselect_n
		.av_ide_read_n       (~mm_interconnect_0_cf_0_ide_read),       //         .read_n
		.av_ide_write_n      (~mm_interconnect_0_cf_0_ide_write),      //         .write_n
		.av_ide_writedata    (mm_interconnect_0_cf_0_ide_writedata),   //         .writedata
		.av_ide_address      (mm_interconnect_0_cf_0_ide_address),     //         .address
		.av_ide_readdata     (mm_interconnect_0_cf_0_ide_readdata),    //         .readdata
		.av_ide_irq          (irq_mapper_receiver1_irq),               //  ide_irq.irq
		.av_ctl_irq          (irq_mapper_receiver0_irq),               //  ctl_irq.irq
		.av_ctl_address      (mm_interconnect_0_cf_0_ctl_address),     //      ctl.address
		.av_ctl_chipselect_n (~mm_interconnect_0_cf_0_ctl_chipselect), //         .chipselect_n
		.av_ctl_read_n       (~mm_interconnect_0_cf_0_ctl_read),       //         .read_n
		.av_ctl_write_n      (~mm_interconnect_0_cf_0_ctl_write),      //         .write_n
		.av_ctl_readdata     (mm_interconnect_0_cf_0_ctl_readdata),    //         .readdata
		.av_ctl_writedata    (mm_interconnect_0_cf_0_ctl_writedata)    //         .writedata
	);

	kernel_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	kernel_epcs epcs (
		.clk           (clk_clk),                                             //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                     //             reset.reset_n
		.reset_req     (rst_controller_reset_out_reset_req),                  //                  .reset_req
		.address       (mm_interconnect_0_epcs_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_0_epcs_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                    //                  .dataavailable
		.endofpacket   (),                                                    //                  .endofpacket
		.read_n        (~mm_interconnect_0_epcs_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_0_epcs_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                    //                  .readyfordata
		.write_n       (~mm_interconnect_0_epcs_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_0_epcs_epcs_control_port_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver4_irq),                            //               irq.irq
		.dclk          (epcs_flash_dclk),                                     //          external.export
		.sce           (epcs_flash_sce),                                      //                  .export
		.sdo           (epcs_flash_sdo),                                      //                  .export
		.data0         (epcs_flash_data0)                                     //                  .export
	);

	kernel_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                   //               irq.irq
	);

	kernel_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	kernel_sdram_ctrl sdram_ctrl (
		.clk            (clk_clk),                                       //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),               // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_ctrl_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_ctrl_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_ctrl_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_ctrl_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_ctrl_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_ctrl_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_ctrl_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_ctrl_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_ctrl_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_ctrl_addr),                               //  wire.export
		.zs_ba          (sdram_ctrl_ba),                                 //      .export
		.zs_cas_n       (sdram_ctrl_cas_n),                              //      .export
		.zs_cke         (sdram_ctrl_cke),                                //      .export
		.zs_cs_n        (sdram_ctrl_cs_n),                               //      .export
		.zs_dq          (sdram_ctrl_dq),                                 //      .export
		.zs_dqm         (sdram_ctrl_dqm),                                //      .export
		.zs_ras_n       (sdram_ctrl_ras_n),                              //      .export
		.zs_we_n        (sdram_ctrl_we_n)                                //      .export
	);

	kernel_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	kernel_uart uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.dataavailable (),                                        //                    .dataavailable
		.readyfordata  (),                                        //                    .readyfordata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver2_irq)                 //                 irq.irq
	);

	kernel_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                             (clk_clk),                                                   //                         clk_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                            // cpu_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                 cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                .readdata
		.cpu_data_master_readdatavalid           (cpu_data_master_readdatavalid),                             //                                .readdatavalid
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //          cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                .readdata
		.cpu_instruction_master_readdatavalid    (cpu_instruction_master_readdatavalid),                      //                                .readdatavalid
		.cf_0_ctl_address                        (mm_interconnect_0_cf_0_ctl_address),                        //                        cf_0_ctl.address
		.cf_0_ctl_write                          (mm_interconnect_0_cf_0_ctl_write),                          //                                .write
		.cf_0_ctl_read                           (mm_interconnect_0_cf_0_ctl_read),                           //                                .read
		.cf_0_ctl_readdata                       (mm_interconnect_0_cf_0_ctl_readdata),                       //                                .readdata
		.cf_0_ctl_writedata                      (mm_interconnect_0_cf_0_ctl_writedata),                      //                                .writedata
		.cf_0_ctl_chipselect                     (mm_interconnect_0_cf_0_ctl_chipselect),                     //                                .chipselect
		.cf_0_ide_address                        (mm_interconnect_0_cf_0_ide_address),                        //                        cf_0_ide.address
		.cf_0_ide_write                          (mm_interconnect_0_cf_0_ide_write),                          //                                .write
		.cf_0_ide_read                           (mm_interconnect_0_cf_0_ide_read),                           //                                .read
		.cf_0_ide_readdata                       (mm_interconnect_0_cf_0_ide_readdata),                       //                                .readdata
		.cf_0_ide_writedata                      (mm_interconnect_0_cf_0_ide_writedata),                      //                                .writedata
		.cf_0_ide_chipselect                     (mm_interconnect_0_cf_0_ide_chipselect),                     //                                .chipselect
		.cpu_debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),             //             cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                .write
		.cpu_debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                .read
		.cpu_debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                .readdata
		.cpu_debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                .writedata
		.cpu_debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                .byteenable
		.cpu_debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                .waitrequest
		.cpu_debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                .debugaccess
		.epcs_epcs_control_port_address          (mm_interconnect_0_epcs_epcs_control_port_address),          //          epcs_epcs_control_port.address
		.epcs_epcs_control_port_write            (mm_interconnect_0_epcs_epcs_control_port_write),            //                                .write
		.epcs_epcs_control_port_read             (mm_interconnect_0_epcs_epcs_control_port_read),             //                                .read
		.epcs_epcs_control_port_readdata         (mm_interconnect_0_epcs_epcs_control_port_readdata),         //                                .readdata
		.epcs_epcs_control_port_writedata        (mm_interconnect_0_epcs_epcs_control_port_writedata),        //                                .writedata
		.epcs_epcs_control_port_chipselect       (mm_interconnect_0_epcs_epcs_control_port_chipselect),       //                                .chipselect
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                .chipselect
		.onchip_memory_s1_address                (mm_interconnect_0_onchip_memory_s1_address),                //                onchip_memory_s1.address
		.onchip_memory_s1_write                  (mm_interconnect_0_onchip_memory_s1_write),                  //                                .write
		.onchip_memory_s1_readdata               (mm_interconnect_0_onchip_memory_s1_readdata),               //                                .readdata
		.onchip_memory_s1_writedata              (mm_interconnect_0_onchip_memory_s1_writedata),              //                                .writedata
		.onchip_memory_s1_byteenable             (mm_interconnect_0_onchip_memory_s1_byteenable),             //                                .byteenable
		.onchip_memory_s1_chipselect             (mm_interconnect_0_onchip_memory_s1_chipselect),             //                                .chipselect
		.onchip_memory_s1_clken                  (mm_interconnect_0_onchip_memory_s1_clken),                  //                                .clken
		.sdram_ctrl_s1_address                   (mm_interconnect_0_sdram_ctrl_s1_address),                   //                   sdram_ctrl_s1.address
		.sdram_ctrl_s1_write                     (mm_interconnect_0_sdram_ctrl_s1_write),                     //                                .write
		.sdram_ctrl_s1_read                      (mm_interconnect_0_sdram_ctrl_s1_read),                      //                                .read
		.sdram_ctrl_s1_readdata                  (mm_interconnect_0_sdram_ctrl_s1_readdata),                  //                                .readdata
		.sdram_ctrl_s1_writedata                 (mm_interconnect_0_sdram_ctrl_s1_writedata),                 //                                .writedata
		.sdram_ctrl_s1_byteenable                (mm_interconnect_0_sdram_ctrl_s1_byteenable),                //                                .byteenable
		.sdram_ctrl_s1_readdatavalid             (mm_interconnect_0_sdram_ctrl_s1_readdatavalid),             //                                .readdatavalid
		.sdram_ctrl_s1_waitrequest               (mm_interconnect_0_sdram_ctrl_s1_waitrequest),               //                                .waitrequest
		.sdram_ctrl_s1_chipselect                (mm_interconnect_0_sdram_ctrl_s1_chipselect),                //                                .chipselect
		.sysid_control_slave_address             (mm_interconnect_0_sysid_control_slave_address),             //             sysid_control_slave.address
		.sysid_control_slave_readdata            (mm_interconnect_0_sysid_control_slave_readdata),            //                                .readdata
		.uart_s1_address                         (mm_interconnect_0_uart_s1_address),                         //                         uart_s1.address
		.uart_s1_write                           (mm_interconnect_0_uart_s1_write),                           //                                .write
		.uart_s1_read                            (mm_interconnect_0_uart_s1_read),                            //                                .read
		.uart_s1_readdata                        (mm_interconnect_0_uart_s1_readdata),                        //                                .readdata
		.uart_s1_writedata                       (mm_interconnect_0_uart_s1_writedata),                       //                                .writedata
		.uart_s1_begintransfer                   (mm_interconnect_0_uart_s1_begintransfer),                   //                                .begintransfer
		.uart_s1_chipselect                      (mm_interconnect_0_uart_s1_chipselect)                       //                                .chipselect
	);

	kernel_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),      // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
